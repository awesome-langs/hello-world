package example where 

example :: Module Empty
example = 
    module 
        let hello =  $display "Hello World!";
        rules 
            "main": when True ==> do 
                hello; 
                $finish 0;